library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
ENTITY dbrom_romonly IS
	port (		addrb: IN std_logic_VECTOR(11 downto 0);
		clkb: IN std_logic;
		dob: OUT std_logic_VECTOR(17 downto 0)	:= (others => '0')
	);
end dbrom_romonly;
architecture behavior of dbrom_romonly is
signal addr : std_logic_vector(11 downto 0):=(others=>'0');
begin
	addr<=addrb;
process(clkb)
begin
	if clkb'event and clkb='1' then
		case addr is
			when "000000000000" => dob<="101010111100010100";
			when "000000000001" => dob<="011100000011110000";
			when "000000000010" => dob<="000001000000000010";
			when "000000000011" => dob<="000110000000000000";
			when "000000000100" => dob<="001001010011011101";
			when "000000000101" => dob<="000000000000000100";
			when "000000000110" => dob<="001110000000010000";
			when "000000000111" => dob<="101010010100010010";
			when "000000001000" => dob<="011100000001010000";
			when "000000001001" => dob<="000110000010101010";
			when "000000001010" => dob<="001001000000001100";
			when "000000001011" => dob<="001000000000100111";
			when "000000001100" => dob<="101010111100010010";
			when "000000001101" => dob<="011100000011110000";
			when "000000001110" => dob<="000110000010101010";
			when "000000001111" => dob<="001001000000010001";
			when "000000010000" => dob<="001000000011011011";
			when "000000010001" => dob<="101010111100010010";
			when "000000010010" => dob<="011100000011110000";
			when "000000010011" => dob<="000110000010101010";
			when "000000010100" => dob<="001001000000010110";
			when "000000010101" => dob<="001000000011011011";
			when "000000010110" => dob<="101010111100010010";
			when "000000010111" => dob<="011100000011110000";
			when "000000011000" => dob<="000110000010101010";
			when "000000011001" => dob<="001001000000011011";
			when "000000011010" => dob<="001000000011011011";
			when "000000011011" => dob<="101010111100010010";
			when "000000011100" => dob<="011100000011110000";
			when "000000011101" => dob<="000110000010101010";
			when "000000011110" => dob<="001001000000100000";
			when "000000011111" => dob<="001000000011011011";
			when "000000100000" => dob<="101010111100010010";
			when "000000100001" => dob<="011100000011110000";
			when "000000100010" => dob<="000110000000000000";
			when "000000100011" => dob<="001001000000100101";
			when "000000100100" => dob<="001000000011011011";
			when "000000100101" => dob<="000000111000000000";
			when "000000100110" => dob<="001000000001101001";
			when "000000100111" => dob<="101010111011111010";
			when "000000101000" => dob<="011100000001010000";
			when "000000101001" => dob<="011100000011100110";
			when "000000101010" => dob<="001001000000101100";
			when "000000101011" => dob<="001000000001001100";
			when "000000101100" => dob<="101010111100010010";
			when "000000101101" => dob<="101010111011111011";
			when "000000101110" => dob<="011100000011110000";
			when "000000101111" => dob<="011100000011100110";
			when "000000110000" => dob<="001001000000110010";
			when "000000110001" => dob<="001000000011011011";
			when "000000110010" => dob<="101010111100010010";
			when "000000110011" => dob<="101010111011111100";
			when "000000110100" => dob<="011100000011110000";
			when "000000110101" => dob<="011100000011100110";
			when "000000110110" => dob<="001001000000111000";
			when "000000110111" => dob<="001000000011011011";
			when "000000111000" => dob<="101010111100010010";
			when "000000111001" => dob<="101010111011111101";
			when "000000111010" => dob<="011100000011110000";
			when "000000111011" => dob<="011100000011100110";
			when "000000111100" => dob<="001001000000111110";
			when "000000111101" => dob<="001000000011011011";
			when "000000111110" => dob<="101010111100010010";
			when "000000111111" => dob<="101010111011111110";
			when "000001000000" => dob<="011100000011110000";
			when "000001000001" => dob<="011100000011100110";
			when "000001000010" => dob<="001001000001000100";
			when "000001000011" => dob<="001000000011011011";
			when "000001000100" => dob<="101010111100010010";
			when "000001000101" => dob<="101010111011111111";
			when "000001000110" => dob<="011100000011110000";
			when "000001000111" => dob<="011100000011100110";
			when "000001001000" => dob<="001001000001001010";
			when "000001001001" => dob<="001000000011011011";
			when "000001001010" => dob<="000000111000000000";
			when "000001001011" => dob<="001000000001101001";
			when "000001001100" => dob<="011100000001010000";
			when "000001001101" => dob<="000110000011111111";
			when "000001001110" => dob<="001001000001010000";
			when "000001001111" => dob<="001000000011011011";
			when "000001010000" => dob<="101010111100010010";
			when "000001010001" => dob<="011100000011110000";
			when "000001010010" => dob<="000110000011111111";
			when "000001010011" => dob<="001001000001010101";
			when "000001010100" => dob<="001000000011011011";
			when "000001010101" => dob<="101010111100010010";
			when "000001010110" => dob<="011100000011110000";
			when "000001010111" => dob<="000110000011111111";
			when "000001011000" => dob<="001001000001011010";
			when "000001011001" => dob<="001000000011011011";
			when "000001011010" => dob<="101010111100010010";
			when "000001011011" => dob<="011100000011110000";
			when "000001011100" => dob<="000110000011111111";
			when "000001011101" => dob<="001001000001011111";
			when "000001011110" => dob<="001000000011011011";
			when "000001011111" => dob<="101010111100010010";
			when "000001100000" => dob<="011100000011110000";
			when "000001100001" => dob<="000110000011111111";
			when "000001100010" => dob<="001001000001100100";
			when "000001100011" => dob<="001000000011011011";
			when "000001100100" => dob<="101010111100010010";
			when "000001100101" => dob<="011100000011110000";
			when "000001100110" => dob<="000110000011111111";
			when "000001100111" => dob<="001001000001101001";
			when "000001101000" => dob<="001000000011011011";
			when "000001101001" => dob<="000000000000010000";
			when "000001101010" => dob<="001110000000010000";
			when "000001101011" => dob<="101010111100010010";
			when "000001101100" => dob<="101010111000010010";
			when "000001101101" => dob<="011100000011110000";
			when "000001101110" => dob<="000110000000001000";
			when "000001101111" => dob<="001001010011011011";
			when "000001110000" => dob<="011100000011100000";
			when "000001110001" => dob<="000110000000001111";
			when "000001110010" => dob<="001001010011011011";
			when "000001110011" => dob<="000000000000010110";
			when "000001110100" => dob<="001110000000010000";
			when "000001110101" => dob<="101010110100010010";
			when "000001110110" => dob<="101010110000010010";
			when "000001110111" => dob<="011100000011000000";
			when "000001111000" => dob<="000110000000000100";
			when "000001111001" => dob<="001001010011011011";
			when "000001111010" => dob<="101010101100010010";
			when "000001111011" => dob<="101010101000010010";
			when "000001111100" => dob<="000000000000011100";
			when "000001111101" => dob<="001110000000010000";
			when "000001111110" => dob<="101010100100010010";
			when "000001111111" => dob<="101010100000010010";
			when "000010000000" => dob<="101110100100100000";
			when "000010000001" => dob<="101110100000100001";
			when "000010000010" => dob<="011100000011010000";
			when "000010000011" => dob<="000110000000000110";
			when "000010000100" => dob<="001001010010001010";
			when "000010000101" => dob<="101010011100010010";
			when "000010000110" => dob<="101010011000010010";
			when "000010000111" => dob<="101110011100100010";
			when "000010001000" => dob<="101110011000100011";
			when "000010001001" => dob<="001000000011011011";
			when "000010001010" => dob<="011100000011010000";
			when "000010001011" => dob<="000110000000000111";
			when "000010001100" => dob<="001001000010010000";
			when "000010001101" => dob<="011100000011010000";
			when "000010001110" => dob<="000110000000001000";
			when "000010001111" => dob<="001001010011011011";
			when "000010010000" => dob<="011100000011010000";
			when "000010010001" => dob<="000110000000000111";
			when "000010010010" => dob<="001001010010010110";
			when "000010010011" => dob<="101010011100100010";
			when "000010010100" => dob<="101010011000100011";
			when "000010010101" => dob<="001000000010011010";
			when "000010010110" => dob<="101010011100010010";
			when "000010010111" => dob<="101010011000010010";
			when "000010011000" => dob<="101110011100100010";
			when "000010011001" => dob<="101110011000100011";
			when "000010011010" => dob<="000000000000000000";
			when "000010011011" => dob<="001110000000000000";
			when "000010011100" => dob<="000000000000111100";
			when "000010011101" => dob<="001110000000000010";
			when "000010011110" => dob<="000000000000111100";
			when "000010011111" => dob<="001110000000000010";
			when "000010100000" => dob<="000000000000000000";
			when "000010100001" => dob<="001110000000000010";
			when "000010100010" => dob<="000000000000000000";
			when "000010100011" => dob<="001110000000000010";
			when "000010100100" => dob<="000000000000000000";
			when "000010100101" => dob<="001110000000000010";
			when "000010100110" => dob<="000000000000000000";
			when "000010100111" => dob<="001110000000000010";
			when "000010101000" => dob<="000000000000000000";
			when "000010101001" => dob<="001110000000000010";
			when "000010101010" => dob<="000000000000000000";
			when "000010101011" => dob<="001110000000000010";
			when "000010101100" => dob<="000000000000001010";
			when "000010101101" => dob<="001110000000010000";
			when "000010101110" => dob<="101010111100010010";
			when "000010101111" => dob<="101110111100000010";
			when "000010110000" => dob<="101010111100010010";
			when "000010110001" => dob<="101110111100000010";
			when "000010110010" => dob<="101010111100010010";
			when "000010110011" => dob<="101110111100000010";
			when "000010110100" => dob<="101010111100010010";
			when "000010110101" => dob<="101110111100000010";
			when "000010110110" => dob<="101010111100010010";
			when "000010110111" => dob<="101110111100000010";
			when "000010111000" => dob<="101010111100010010";
			when "000010111001" => dob<="101110111100000010";
			when "000010111010" => dob<="000000000010101010";
			when "000010111011" => dob<="001110000000000010";
			when "000010111100" => dob<="000000000010101010";
			when "000010111101" => dob<="001110000000000010";
			when "000010111110" => dob<="000000000010101010";
			when "000010111111" => dob<="001110000000000010";
			when "000011000000" => dob<="000000000010101010";
			when "000011000001" => dob<="001110000000000010";
			when "000011000010" => dob<="000000000010101010";
			when "000011000011" => dob<="001110000000000010";
			when "000011000100" => dob<="000000000000000000";
			when "000011000101" => dob<="001110000000000010";
			when "000011000110" => dob<="000000000000001000";
			when "000011000111" => dob<="001110000000000010";
			when "000011001000" => dob<="000000000000001011";
			when "000011001001" => dob<="001110000000000010";
			when "000011001010" => dob<="000000000000011010";
			when "000011001011" => dob<="001110000000000000";
			when "000011001100" => dob<="101110110100000010";
			when "000011001101" => dob<="000000000010000100";
			when "000011001110" => dob<="001110000000000010";
			when "000011001111" => dob<="101110101100000010";
			when "000011010000" => dob<="101110101000000010";
			when "000011010001" => dob<="000000000000000100";
			when "000011010010" => dob<="001110000000000010";
			when "000011010011" => dob<="000000000000000000";
			when "000011010100" => dob<="001110000000000010";
			when "000011010101" => dob<="101110100100000010";
			when "000011010110" => dob<="101110100000000010";
			when "000011010111" => dob<="101110011100000010";
			when "000011011000" => dob<="101110011000000010";
			when "000011011001" => dob<="000000000000000000";
			when "000011011010" => dob<="001110000000001000";
			when "000011011011" => dob<="000000000000000000";
			when "000011011100" => dob<="001110000000011010";
			when "000011011101" => dob<="001000000000000000";
			when "000011011110" => dob<="001000100000000000";
			when others => dob<="000000000000000000";
		end case;
	end if;
end process;
end behavior;
