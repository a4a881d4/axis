library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
ENTITY ethrxrom_romonly IS
	port (		addrb: IN std_logic_VECTOR(11 downto 0);
		clkb: IN std_logic;
		dob: OUT std_logic_VECTOR(17 downto 0)	:= (others => '0')
	);
end ethrxrom_romonly;
architecture behavior of ethrxrom_romonly is
signal addr : std_logic_vector(11 downto 0):=(others=>'0');
begin
	addr<=addrb;
process(clkb)
begin
	if clkb'event and clkb='1' then
		case addr is
			when "000000000000" => dob<="001000110000000100";
			when "000000000001" => dob<="001000110000010110";
			when "000000000010" => dob<="001000000000000001";
			when "000000000011" => dob<="001000100000000000";
			when "000000000100" => dob<="000000000000000000";
			when "000000000101" => dob<="001110000000100011";
			when "000000000110" => dob<="000000000000000000";
			when "000000000111" => dob<="001110000000100100";
			when "000000001000" => dob<="000000000000000000";
			when "000000001001" => dob<="001110000000100101";
			when "000000001010" => dob<="000000000000000000";
			when "000000001011" => dob<="001110000000100111";
			when "000000001100" => dob<="000000000000000000";
			when "000000001101" => dob<="001110000000101000";
			when "000000001110" => dob<="000000000000000000";
			when "000000001111" => dob<="001110000000101001";
			when "000000010000" => dob<="000000000000000001";
			when "000000010001" => dob<="001110000000101011";
			when "000000010010" => dob<="000000000000000001";
			when "000000010011" => dob<="001110000000101100";
			when "000000010100" => dob<="100000010100000000";
			when "000000010101" => dob<="001000100000000000";
			when "000000010110" => dob<="101010111100010100";
			when "000000010111" => dob<="011100000011110000";
			when "000000011000" => dob<="000001000000000010";
			when "000000011001" => dob<="000110000000000000";
			when "000000011010" => dob<="001001010100011100";
			when "000000011011" => dob<="000000000000000100";
			when "000000011100" => dob<="001110000000010000";
			when "000000011101" => dob<="101010000000010010";
			when "000000011110" => dob<="101010111011111001";
			when "000000011111" => dob<="011100000000000000";
			when "000000100000" => dob<="011100000011100110";
			when "000000100001" => dob<="001001000000100011";
			when "000000100010" => dob<="001000000001000010";
			when "000000100011" => dob<="101010111100010010";
			when "000000100100" => dob<="101010111011111011";
			when "000000100101" => dob<="011100000011110000";
			when "000000100110" => dob<="011100000011100110";
			when "000000100111" => dob<="001001000000101001";
			when "000000101000" => dob<="001000000100011010";
			when "000000101001" => dob<="101010111100010010";
			when "000000101010" => dob<="101010111011111100";
			when "000000101011" => dob<="011100000011110000";
			when "000000101100" => dob<="011100000011100110";
			when "000000101101" => dob<="001001000000101111";
			when "000000101110" => dob<="001000000100011010";
			when "000000101111" => dob<="101010111100010010";
			when "000000110000" => dob<="101010111011111101";
			when "000000110001" => dob<="011100000011110000";
			when "000000110010" => dob<="011100000011100110";
			when "000000110011" => dob<="001001000000110101";
			when "000000110100" => dob<="001000000100011010";
			when "000000110101" => dob<="101010111100010010";
			when "000000110110" => dob<="101010111011111110";
			when "000000110111" => dob<="011100000011110000";
			when "000000111000" => dob<="011100000011100110";
			when "000000111001" => dob<="001001000000111011";
			when "000000111010" => dob<="001000000100011010";
			when "000000111011" => dob<="101010111100010010";
			when "000000111100" => dob<="101010111011111111";
			when "000000111101" => dob<="011100000011110000";
			when "000000111110" => dob<="011100000011100110";
			when "000000111111" => dob<="001001000001000001";
			when "000001000000" => dob<="001000000100011010";
			when "000001000001" => dob<="001000000010000011";
			when "000001000010" => dob<="101010111011111010";
			when "000001000011" => dob<="011100000000000000";
			when "000001000100" => dob<="011100000011100110";
			when "000001000101" => dob<="001001000001000111";
			when "000001000110" => dob<="001000000001100110";
			when "000001000111" => dob<="101010111100010010";
			when "000001001000" => dob<="101010111011111011";
			when "000001001001" => dob<="011100000011110000";
			when "000001001010" => dob<="011100000011100110";
			when "000001001011" => dob<="001001000001001101";
			when "000001001100" => dob<="001000000100011010";
			when "000001001101" => dob<="101010111100010010";
			when "000001001110" => dob<="101010111011111100";
			when "000001001111" => dob<="011100000011110000";
			when "000001010000" => dob<="011100000011100110";
			when "000001010001" => dob<="001001000001010011";
			when "000001010010" => dob<="001000000100011010";
			when "000001010011" => dob<="101010111100010010";
			when "000001010100" => dob<="101010111011111101";
			when "000001010101" => dob<="011100000011110000";
			when "000001010110" => dob<="011100000011100110";
			when "000001010111" => dob<="001001000001011001";
			when "000001011000" => dob<="001000000100011010";
			when "000001011001" => dob<="101010111100010010";
			when "000001011010" => dob<="101010111011111110";
			when "000001011011" => dob<="011100000011110000";
			when "000001011100" => dob<="011100000011100110";
			when "000001011101" => dob<="001001000001011111";
			when "000001011110" => dob<="001000000100011010";
			when "000001011111" => dob<="101010111100010010";
			when "000001100000" => dob<="101010111011111111";
			when "000001100001" => dob<="011100000011110000";
			when "000001100010" => dob<="011100000011100110";
			when "000001100011" => dob<="001001000001100101";
			when "000001100100" => dob<="001000000100011010";
			when "000001100101" => dob<="001000000010000011";
			when "000001100110" => dob<="011100000000000000";
			when "000001100111" => dob<="000110000011111111";
			when "000001101000" => dob<="001001000001101010";
			when "000001101001" => dob<="001000000100011010";
			when "000001101010" => dob<="101010111100010010";
			when "000001101011" => dob<="011100000011110000";
			when "000001101100" => dob<="000110000011111111";
			when "000001101101" => dob<="001001000001101111";
			when "000001101110" => dob<="001000000100011010";
			when "000001101111" => dob<="101010111100010010";
			when "000001110000" => dob<="011100000011110000";
			when "000001110001" => dob<="000110000011111111";
			when "000001110010" => dob<="001001000001110100";
			when "000001110011" => dob<="001000000100011010";
			when "000001110100" => dob<="101010111100010010";
			when "000001110101" => dob<="011100000011110000";
			when "000001110110" => dob<="000110000011111111";
			when "000001110111" => dob<="001001000001111001";
			when "000001111000" => dob<="001000000100011010";
			when "000001111001" => dob<="101010111100010010";
			when "000001111010" => dob<="011100000011110000";
			when "000001111011" => dob<="000110000011111111";
			when "000001111100" => dob<="001001000001111110";
			when "000001111101" => dob<="001000000100011010";
			when "000001111110" => dob<="101010111100010010";
			when "000001111111" => dob<="011100000011110000";
			when "000010000000" => dob<="000110000011111111";
			when "000010000001" => dob<="001001000010000011";
			when "000010000010" => dob<="001000000100011010";
			when "000010000011" => dob<="000000000000010000";
			when "000010000100" => dob<="001110000000010000";
			when "000010000101" => dob<="101010111000010010";
			when "000010000110" => dob<="101010111100010010";
			when "000010000111" => dob<="011100000011100000";
			when "000010001000" => dob<="000110000000001000";
			when "000010001001" => dob<="001001010011011100";
			when "000010001010" => dob<="011100000011110000";
			when "000010001011" => dob<="000110000000001010";
			when "000010001100" => dob<="001001010011011100";
			when "000010001101" => dob<="000000000000010110";
			when "000010001110" => dob<="001110000000010000";
			when "000010001111" => dob<="101010110100010010";
			when "000010010000" => dob<="101010101000010010";
			when "000010010001" => dob<="101010100100010010";
			when "000010010010" => dob<="101010100000010010";
			when "000010010011" => dob<="101010011100010010";
			when "000010010100" => dob<="101110101000100111";
			when "000010010101" => dob<="101110100100101000";
			when "000010010110" => dob<="101110100000101001";
			when "000010010111" => dob<="101110011100101010";
			when "000010011000" => dob<="011100000011010000";
			when "000010011001" => dob<="000001000000000001";
			when "000010011010" => dob<="000110000000000000";
			when "000010011011" => dob<="001001000010101111";
			when "000010011100" => dob<="000000000000011111";
			when "000010011101" => dob<="001110000000010000";
			when "000010011110" => dob<="101010111100010010";
			when "000010011111" => dob<="000000000000000000";
			when "000010100000" => dob<="011100000011110110";
			when "000010100001" => dob<="001001110010100101";
			when "000010100010" => dob<="111100110011110000";
			when "000010100011" => dob<="100000101100000000";
			when "000010100100" => dob<="001000000010101110";
			when "000010100101" => dob<="000000000000000000";
			when "000010100110" => dob<="001110000000010000";
			when "000010100111" => dob<="101010110000010010";
			when "000010101000" => dob<="101010101100010010";
			when "000010101001" => dob<="011100000011000000";
			when "000010101010" => dob<="000110000000100100";
			when "000010101011" => dob<="001001110010101101";
			when "000010101100" => dob<="100110101100000001";
			when "000010101101" => dob<="100110110000100100";
			when "000010101110" => dob<="001000000010111000";
			when "000010101111" => dob<="000000000000000000";
			when "000010110000" => dob<="001110000000010000";
			when "000010110001" => dob<="101010110000010010";
			when "000010110010" => dob<="101010101100010010";
			when "000010110011" => dob<="011100000011000000";
			when "000010110100" => dob<="000110000000011000";
			when "000010110101" => dob<="001001110010110111";
			when "000010110110" => dob<="100110101100000001";
			when "000010110111" => dob<="100110110000011000";
			when "000010111000" => dob<="101110110000100001";
			when "000010111001" => dob<="101110101100100010";
			when "000010111010" => dob<="000000000000000010";
			when "000010111011" => dob<="001110000000010000";
			when "000010111100" => dob<="101010111100010010";
			when "000010111101" => dob<="101010111000010010";
			when "000010111110" => dob<="011100000011010000";
			when "000010111111" => dob<="000001000000000001";
			when "000011000000" => dob<="000110000000000000";
			when "000011000001" => dob<="001001000011001000";
			when "000011000010" => dob<="100100111100100100";
			when "000011000011" => dob<="011100000011110000";
			when "000011000100" => dob<="000110000000100100";
			when "000011000101" => dob<="001001110011000111";
			when "000011000110" => dob<="100100111000000001";
			when "000011000111" => dob<="001000000011001101";
			when "000011001000" => dob<="100100111100011000";
			when "000011001001" => dob<="011100000011110000";
			when "000011001010" => dob<="000110000000011000";
			when "000011001011" => dob<="001001110011001101";
			when "000011001100" => dob<="100100111000000001";
			when "000011001101" => dob<="101110111100100011";
			when "000011001110" => dob<="101110111000100100";
			when "000011001111" => dob<="101010111000101101";
			when "000011010000" => dob<="011100000011100000";
			when "000011010001" => dob<="000001000000000001";
			when "000011010010" => dob<="000110000000000000";
			when "000011010011" => dob<="001001010011001111";
			when "000011010100" => dob<="000000000000000000";
			when "000011010101" => dob<="001110000000100000";
			when "000011010110" => dob<="011100000011010000";
			when "000011010111" => dob<="000001000000000001";
			when "000011011000" => dob<="000110000000000000";
			when "000011011001" => dob<="001001000011011011";
			when "000011011010" => dob<="001000110100011101";
			when "000011011011" => dob<="001000000100011010";
			when "000011011100" => dob<="011100000011100000";
			when "000011011101" => dob<="000110000000001000";
			when "000011011110" => dob<="001001010100011010";
			when "000011011111" => dob<="011100000011110000";
			when "000011100000" => dob<="000110000000001011";
			when "000011100001" => dob<="001001010100011010";
			when "000011100010" => dob<="101010111100110100";
			when "000011100011" => dob<="011100000011110000";
			when "000011100100" => dob<="000001000000000001";
			when "000011100101" => dob<="000110000000000000";
			when "000011100110" => dob<="001001010011100010";
			when "000011100111" => dob<="000000000000011100";
			when "000011101000" => dob<="001110000000010000";
			when "000011101001" => dob<="101010111100010010";
			when "000011101010" => dob<="101010111000010010";
			when "000011101011" => dob<="000000000000000000";
			when "000011101100" => dob<="001110000000110000";
			when "000011101101" => dob<="101110111100110010";
			when "000011101110" => dob<="101110111000110010";
			when "000011101111" => dob<="101010111100010010";
			when "000011110000" => dob<="101010111000010010";
			when "000011110001" => dob<="101110111100110010";
			when "000011110010" => dob<="101110111000110010";
			when "000011110011" => dob<="000000000000010110";
			when "000011110100" => dob<="001110000000010000";
			when "000011110101" => dob<="101010111100010010";
			when "000011110110" => dob<="000000000000000000";
			when "000011110111" => dob<="001110000000110010";
			when "000011111000" => dob<="000000000000000000";
			when "000011111001" => dob<="001110000000110010";
			when "000011111010" => dob<="000000000000000000";
			when "000011111011" => dob<="001110000000110010";
			when "000011111100" => dob<="011100000011110000";
			when "000011111101" => dob<="000110000000000110";
			when "000011111110" => dob<="001001010100000010";
			when "000011111111" => dob<="000000000000000000";
			when "000100000000" => dob<="001110000000110010";
			when "000100000001" => dob<="001000000100000111";
			when "000100000010" => dob<="011100000011110000";
			when "000100000011" => dob<="000110000000000111";
			when "000100000100" => dob<="001001010100000111";
			when "000100000101" => dob<="000000000000000001";
			when "000100000110" => dob<="001110000000110010";
			when "000100000111" => dob<="000000000000001100";
			when "000100001000" => dob<="001110000000110000";
			when "000100001001" => dob<="000000000000001010";
			when "000100001010" => dob<="001110000000010000";
			when "000100001011" => dob<="101010011000010010";
			when "000100001100" => dob<="101110011000110010";
			when "000100001101" => dob<="101010011000010010";
			when "000100001110" => dob<="101110011000110010";
			when "000100001111" => dob<="101010011000010010";
			when "000100010000" => dob<="101110011000110010";
			when "000100010001" => dob<="101010011000010010";
			when "000100010010" => dob<="101110011000110010";
			when "000100010011" => dob<="101010011000010010";
			when "000100010100" => dob<="101110011000110010";
			when "000100010101" => dob<="101010011000010010";
			when "000100010110" => dob<="101110011000110010";
			when "000100010111" => dob<="101110000000110010";
			when "000100011000" => dob<="000000000000000000";
			when "000100011001" => dob<="001110000000111000";
			when "000100011010" => dob<="000000000000000000";
			when "000100011011" => dob<="001110000000011010";
			when "000100011100" => dob<="001000100000000000";
			when "000100011101" => dob<="101010111100110100";
			when "000100011110" => dob<="011100000011110000";
			when "000100011111" => dob<="000001000000000001";
			when "000100100000" => dob<="000110000000000000";
			when "000100100001" => dob<="001001010100011101";
			when "000100100010" => dob<="000000000000100000";
			when "000100100011" => dob<="001110000000010000";
			when "000100100100" => dob<="101010101000010010";
			when "000100100101" => dob<="101010100100010010";
			when "000100100110" => dob<="101010100000010010";
			when "000100100111" => dob<="101010011100010010";
			when "000100101000" => dob<="000000000000000000";
			when "000100101001" => dob<="001110000000110000";
			when "000100101010" => dob<="101110011100110010";
			when "000100101011" => dob<="101110100000110010";
			when "000100101100" => dob<="101110100100110010";
			when "000100101101" => dob<="101110101000110010";
			when "000100101110" => dob<="101010010000010010";
			when "000100101111" => dob<="101010001100010010";
			when "000100110000" => dob<="101010001000010010";
			when "000100110001" => dob<="101010000100010010";
			when "000100110010" => dob<="101110000100110010";
			when "000100110011" => dob<="101110001000110010";
			when "000100110100" => dob<="101110001100110010";
			when "000100110101" => dob<="101110010000110010";
			when "000100110110" => dob<="000000000000011011";
			when "000100110111" => dob<="001110000000010000";
			when "000100111000" => dob<="101010011000010010";
			when "000100111001" => dob<="101110011000110010";
			when "000100111010" => dob<="101010011000010010";
			when "000100111011" => dob<="101110011000110010";
			when "000100111100" => dob<="101010011000010010";
			when "000100111101" => dob<="101110011000110010";
			when "000100111110" => dob<="101010011000010010";
			when "000100111111" => dob<="101110011000110010";
			when "000101000000" => dob<="000000000000001010";
			when "000101000001" => dob<="001110000000010000";
			when "000101000010" => dob<="101010011000010010";
			when "000101000011" => dob<="101110011000110010";
			when "000101000100" => dob<="101010011000010010";
			when "000101000101" => dob<="101110011000110010";
			when "000101000110" => dob<="101010011000010010";
			when "000101000111" => dob<="101110011000110010";
			when "000101001000" => dob<="101010011000010010";
			when "000101001001" => dob<="101110011000110010";
			when "000101001010" => dob<="101010011000010010";
			when "000101001011" => dob<="101110011000110010";
			when "000101001100" => dob<="101010011000010010";
			when "000101001101" => dob<="101110011000110010";
			when "000101001110" => dob<="101110000000110010";
			when "000101001111" => dob<="000000000000000000";
			when "000101010000" => dob<="001110000000101110";
			when "000101010001" => dob<="100000010100000000";
			when "000101010010" => dob<="001000100000000000";
			when others => dob<="000000000000000000";
		end case;
	end if;
end process;
end behavior;
